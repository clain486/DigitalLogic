module alu(a,b,aluc,r,zero,carry,negative,overflow);
input [31:0] a,b;
input [3:0] aluc;
output reg [31:0] r;
output reg zero,carry,negative,overflow;

always@(*)
begin
    case(aluc)
        //add
        4'b0010:
            begin
            r=a+b;
            overflow=((a[31]==b[31])&&(~r[31]==a[31]))?1:0;
            zero=(r==0)?1:0;
            carry=0;
            negative=(r<0)?1:0;
            end
        //addu
        4'b0000:
            begin
            {carry,r}=a+b;
            zero=(r==0)?1:0;
            overflow=0;
            negative=(r[31]==1)?1:0;
            end
        //sub
        4'b0011:
            begin
            r=a-b;
            overflow=((a[31]==0 && b[31]==1 && r[31]==1) || (a[31]==1 && b[31]==0 && r[31]==0))?1:0;
            zero=(a==b)?1:0;
            carry=0;
            negative=(r<0)?1:0;
            end
        //subu
        4'b0001:
            begin
            {carry,r}=a-b;
            zero=(r==0)?1:0;
            overflow=0;
            negative=(r[31]==1)?1:0;
            end
        //and
        4'b0100:
            begin
            r=a&b;
            zero=(r==0)?1:0;
            carry=0;
            overflow=0;
            negative=(r[31]==1)?1:0;
            end
        //or
        4'b0101:
            begin
            r=a|b;
            zero=(r==0)?1:0;
            carry=0;
            overflow=0;
            negative=(r[31]==1)?1:0;
            end
        //xor
        4'b0110:
            begin
            r=a^b;
            zero=(r==0)?1:0;
            carry=0;
            overflow=0;
            negative=(r[31]==1)?1:0;
            end
        //nor
        4'b0111:
            begin
            r=~(a|b);
            zero=(r==0)?1:0;
            carry=0;
            overflow=0;
            negative=(r[31]==1)?1:0;
            end
        //slt
        11'b1011:
            begin                        
            if(a[31]==1 && b[31]==0)
                r=1;
            else if(a[31]==0 && b[31]==1)
                r=0;
            else 
                r=(a<b)?1:0;
           overflow=r; 
           zero=(r==0)?1:0;
           carry=0;
           negative=(a<b)?1:0;
           end
        //sltu
        4'b1010:
            begin
            r=(a<b)?1:0;
            carry=r;
            zero=(r==0)?1:0;
            overflow=0;
            negative=(r[31]==1)?1:0;
            end
        //sll/slr
        4'b111x:
            begin
            {carry,r}=b<<a;
            overflow=0;
            zero=(r==0)?1:0;
            negative=(r[31]==1)?1:0;
            end
        //srl
        4'b1101:
            begin
            r=b>>a;
            carry=b[a-1];
            overflow=0;
            zero=(r==0)?1:0;
            negative=(r[31]==1)?1:0;
            end
        //sra
        4'b1100:
            begin
            r=($signed(b))>>>a;
            carry=b[a];
            overflow=0;
            zero=(r==0)?1:0;
            negative=(r[31]==1)?1:0;
            end
        //lui
        4'b100x:
            begin
            r={b[15:0],16'b0};
            carry=0;
            overflow=0;
            zero=(r==0)?1:0;
            negative=(r[31]==1)?1:0;
            end       
    endcase
end
endmodule
